/*Note:
Mesh input B connected PE input D. Therefore, in mesh B is 16 bits.
Mesh input D connected PE input B. Therefore, in mesh D is 8 bits.
*/

module Mesh( 
  input         clock, 
  //input A, one for each column
  input  [7:0]  io_in_a_0_0, 
  input  [7:0]  io_in_a_1_0, 
  input  [7:0]  io_in_a_2_0, 
  input  [7:0]  io_in_a_3_0, 
  //input B, one for each row
  input  [7:0]  io_in_d_0_0, 
  input  [7:0]  io_in_d_1_0, 
  input  [7:0]  io_in_d_2_0, 
  input  [7:0]  io_in_d_3_0, 
  //input D, for taking output 
  input  [15:0]  io_in_b_0_0, 
  input  [15:0]  io_in_b_1_0, 
  input  [15:0]  io_in_b_2_0, 
  input  [15:0]  io_in_b_3_0, 
  //CTL_PROP, one for each column
  input         io_in_control_0_0_propagate, 
  input         io_in_control_1_0_propagate, 
  input         io_in_control_2_0_propagate, 
  input         io_in_control_3_0_propagate, 
  //Ouputs C_OUT, one from each column at bottom
  output reg [15:0] io_out_c_0_0, 
  output reg [15:0] io_out_c_1_0, 
  output reg [15:0] io_out_c_2_0, 
  output reg [15:0] io_out_c_3_0
 );
 
 //Mesh Internal input/ouput wires intialization
  wire  mesh_0_0_clock; 		  			
  wire [7:0] mesh_0_0_io_in_a_0;  			
  wire [7:0] mesh_0_0_io_in_b_0; 			
  wire [15:0] mesh_0_0_io_in_d_0; 			
  wire  mesh_0_0_io_in_control_0_propagate; 
  wire [7:0] mesh_0_0_io_out_a_0; 			
  wire [15:0] mesh_0_0_io_out_c_0;			
  wire [7:0] mesh_0_0_io_out_b_0;			
  wire  mesh_0_0_io_out_control_0_propagate;
  wire  mesh_0_1_clock; 
  wire [7:0] mesh_0_1_io_in_a_0; 
  wire [7:0] mesh_0_1_io_in_b_0;
  wire [15:0] mesh_0_1_io_in_d_0;
  wire  mesh_0_1_io_in_control_0_propagate; 
  wire [7:0] mesh_0_1_io_out_a_0; 
  wire [15:0] mesh_0_1_io_out_c_0;
  wire [7:0] mesh_0_1_io_out_b_0;
  wire  mesh_0_1_io_out_control_0_propagate; 
  wire  mesh_0_2_clock; 			
  wire [7:0] mesh_0_2_io_in_a_0; 	
  wire [7:0] mesh_0_2_io_in_b_0; 	
  wire [15:0] mesh_0_2_io_in_d_0; 	
  wire  mesh_0_2_io_in_control_0_propagate; 
  wire [7:0] mesh_0_2_io_out_a_0; 
  wire [15:0] mesh_0_2_io_out_c_0;
  wire [7:0] mesh_0_2_io_out_b_0;
  wire  mesh_0_2_io_out_control_0_propagate; 
  wire  mesh_0_3_clock; 		 
  wire [7:0] mesh_0_3_io_in_a_0; 
  wire [7:0] mesh_0_3_io_in_b_0;
  wire [15:0] mesh_0_3_io_in_d_0;
  wire  mesh_0_3_io_in_control_0_propagate; 
  wire [7:0] mesh_0_3_io_out_a_0; 
  wire [15:0] mesh_0_3_io_out_c_0;
  wire [7:0] mesh_0_3_io_out_b_0;
  wire  mesh_0_3_io_out_control_0_propagate; 
  
  wire  mesh_1_0_clock;
  wire [7:0] mesh_1_0_io_in_a_0; 
  wire [7:0] mesh_1_0_io_in_b_0;
  wire [15:0] mesh_1_0_io_in_d_0;
  wire  mesh_1_0_io_in_control_0_propagate; 
  wire [7:0] mesh_1_0_io_out_a_0; 
  wire [15:0] mesh_1_0_io_out_c_0;
  wire [7:0] mesh_1_0_io_out_b_0;
  wire  mesh_1_0_io_out_control_0_propagate;
  wire  mesh_1_1_clock; 		 
  wire [7:0] mesh_1_1_io_in_a_0; 
  wire [7:0] mesh_1_1_io_in_b_0;
  wire [15:0] mesh_1_1_io_in_d_0;
  wire  mesh_1_1_io_in_control_0_propagate; 
  wire [7:0] mesh_1_1_io_out_a_0; 			
  wire [15:0] mesh_1_1_io_out_c_0;			
  wire [7:0] mesh_1_1_io_out_b_0;			
  wire  mesh_1_1_io_out_control_0_propagate;
  wire  mesh_1_2_clock; 
  wire [7:0] mesh_1_2_io_in_a_0; 
  wire [7:0] mesh_1_2_io_in_b_0;
  wire [15:0] mesh_1_2_io_in_d_0;
  wire  mesh_1_2_io_in_control_0_propagate; 
  wire [7:0] mesh_1_2_io_out_a_0; 
  wire [15:0] mesh_1_2_io_out_c_0;
  wire [7:0] mesh_1_2_io_out_b_0;
  wire  mesh_1_2_io_out_control_0_propagate;
  wire  mesh_1_3_clock; 		 
  wire [7:0] mesh_1_3_io_in_a_0; 
  wire [7:0] mesh_1_3_io_in_b_0;
  wire [15:0] mesh_1_3_io_in_d_0;
  wire  mesh_1_3_io_in_control_0_propagate; 
  wire [7:0] mesh_1_3_io_out_a_0; 
  wire [15:0] mesh_1_3_io_out_c_0;
  wire [7:0] mesh_1_3_io_out_b_0;
  wire  mesh_1_3_io_out_control_0_propagate;
  
  wire  mesh_2_0_clock; 
  wire [7:0] mesh_2_0_io_in_a_0; 
  wire [7:0] mesh_2_0_io_in_b_0;
  wire [15:0] mesh_2_0_io_in_d_0;
  wire  mesh_2_0_io_in_control_0_propagate; 
  wire [7:0] mesh_2_0_io_out_a_0; 			
  wire [15:0] mesh_2_0_io_out_c_0;			
  wire [7:0] mesh_2_0_io_out_b_0;			
  wire  mesh_2_0_io_out_control_0_propagate;
  wire  mesh_2_1_clock;						
  wire [7:0] mesh_2_1_io_in_a_0; 			
  wire [7:0] mesh_2_1_io_in_b_0;			
  wire [15:0] mesh_2_1_io_in_d_0;			
  wire  mesh_2_1_io_in_control_0_propagate; 
  wire [7:0] mesh_2_1_io_out_a_0; 			
  wire [15:0] mesh_2_1_io_out_c_0;			
  wire [7:0] mesh_2_1_io_out_b_0;			
  wire  mesh_2_1_io_out_control_0_propagate;
  wire  mesh_2_2_clock; 		 			
  wire [7:0] mesh_2_2_io_in_a_0; 			
  wire [7:0] mesh_2_2_io_in_b_0;			
  wire [15:0] mesh_2_2_io_in_d_0;			
  wire  mesh_2_2_io_in_control_0_propagate; 
  wire [7:0] mesh_2_2_io_out_a_0; 			
  wire [15:0] mesh_2_2_io_out_c_0;			
  wire [7:0] mesh_2_2_io_out_b_0;			
  wire  mesh_2_2_io_out_control_0_propagate;
  wire  mesh_2_3_clock; 		 			
  wire [7:0] mesh_2_3_io_in_a_0; 			
  wire [7:0] mesh_2_3_io_in_b_0;			
  wire [15:0] mesh_2_3_io_in_d_0;			
  wire  mesh_2_3_io_in_control_0_propagate; 
  wire [7:0] mesh_2_3_io_out_a_0; 			
  wire [15:0] mesh_2_3_io_out_c_0;			
  wire [7:0] mesh_2_3_io_out_b_0;			
  wire  mesh_2_3_io_out_control_0_propagate;
  
  wire  mesh_3_0_clock;			 
  wire [7:0] mesh_3_0_io_in_a_0; 
  wire [7:0] mesh_3_0_io_in_b_0;
  wire [15:0] mesh_3_0_io_in_d_0;
  wire  mesh_3_0_io_in_control_0_propagate; 
  wire [7:0] mesh_3_0_io_out_a_0; 
  wire [15:0] mesh_3_0_io_out_c_0;
  wire [7:0] mesh_3_0_io_out_b_0;
  wire  mesh_3_0_io_out_control_0_propagate;
  wire  mesh_3_1_clock; 		 
  wire [7:0] mesh_3_1_io_in_a_0; 
  wire [7:0] mesh_3_1_io_in_b_0;
  wire [15:0] mesh_3_1_io_in_d_0;
  wire  mesh_3_1_io_in_control_0_propagate; 
  wire [7:0] mesh_3_1_io_out_a_0; 
  wire [15:0] mesh_3_1_io_out_c_0;
  wire [7:0] mesh_3_1_io_out_b_0;
  wire  mesh_3_1_io_out_control_0_propagate;
  wire  mesh_3_2_clock; 
  wire [7:0] mesh_3_2_io_in_a_0; 
  wire [7:0] mesh_3_2_io_in_b_0;
  wire [15:0] mesh_3_2_io_in_d_0;
  wire  mesh_3_2_io_in_control_0_propagate; 
  wire [7:0] mesh_3_2_io_out_a_0; 
  wire [15:0] mesh_3_2_io_out_c_0;
  wire [7:0] mesh_3_2_io_out_b_0;
  wire  mesh_3_2_io_out_control_0_propagate;
  wire  mesh_3_3_clock;
  wire [7:0] mesh_3_3_io_in_a_0; 
  wire [7:0] mesh_3_3_io_in_b_0;
  wire [15:0] mesh_3_3_io_in_d_0;
  wire  mesh_3_3_io_in_control_0_propagate; 
  wire [7:0] mesh_3_3_io_out_a_0; 
  wire [15:0] mesh_3_3_io_out_c_0;
  wire [7:0] mesh_3_3_io_out_b_0;
  wire  mesh_3_3_io_out_control_0_propagate;
  

//I/O Registers initialization 
  reg [7:0] _T_1_0; 
  reg [31:0] _RAND_1;
  reg [7:0] _T_2_0; 
  reg [31:0] _RAND_2;
  reg [7:0] _T_3_0; 
  reg [31:0] _RAND_3;
  reg [7:0] _T_4_0; 
  reg [31:0] _RAND_4;

  reg [7:0] _T_10_0;
  reg [31:0] _RAND_10;
  reg [7:0] _T_11_0;
  reg [31:0] _RAND_11;
  reg [7:0] _T_12_0; 
  reg [31:0] _RAND_12;
  reg [7:0] _T_13_0; 
  reg [31:0] _RAND_13;

  reg [7:0] _T_19_0; 
  reg [31:0] _RAND_19;
  reg [7:0] _T_20_0; 
  reg [31:0] _RAND_20;
  reg [7:0] _T_21_0; 
  reg [31:0] _RAND_21;
  reg [7:0] _T_22_0; 
  reg [31:0] _RAND_22;

  reg [7:0] _T_28_0;  
  reg [31:0] _RAND_28;
  reg [7:0] _T_29_0;  
  reg [31:0] _RAND_29;
  reg [7:0] _T_30_0;  
  reg [31:0] _RAND_30;
  reg [7:0] _T_31_0;  
  reg [31:0] _RAND_31;
  
  

  reg [7:0]  _T_74_0;
  reg [31:0] _RAND_74;
  reg [7:0]  _T_75_0; 
  reg [31:0] _RAND_75;
  reg [7:0]  _T_76_0; 
  reg [31:0] _RAND_76;
  reg [7:0]  _T_77_0; 
  reg [31:0] _RAND_77;

  reg [7:0]  _T_84_0;
  reg [31:0] _RAND_84;
  reg [7:0]  _T_85_0; 
  reg [31:0] _RAND_85;
  reg [7:0]  _T_86_0; 
  reg [31:0] _RAND_86;
  reg [7:0]  _T_87_0; 
  reg [31:0] _RAND_87;

  reg [7:0]  _T_94_0; 
  reg [31:0] _RAND_94;
  reg [7:0]  _T_95_0; 
  reg [31:0] _RAND_95;
  reg [7:0]  _T_96_0; 
  reg [31:0] _RAND_96;
  reg [7:0]  _T_97_0; 
  reg [31:0] _RAND_97;
  reg [7:0]  _T_98_0; 
  reg [31:0] _RAND_98;
  reg [7:0]  _T_99_0; 
  reg [31:0] _RAND_99;
  reg [7:0]  _T_100_0;
  reg [31:0] _RAND_100;
  reg [7:0]  _T_101_0; 
  reg [31:0] _RAND_101;

  reg [7:0]  _T_104_0; 
  reg [31:0] _RAND_104;
  reg [7:0]  _T_105_0; 
  reg [31:0] _RAND_105;
  reg [7:0]  _T_106_0; 
  reg [31:0] _RAND_106;
  reg [7:0]  _T_107_0; 
  reg [31:0] _RAND_107;
  

  reg [15:0] _T_154_0;
  reg [31:0] _RAND_154;
  reg [15:0] _T_155_0; 
  reg [31:0] _RAND_155;
  reg [15:0] _T_156_0; 
  reg [31:0] _RAND_156;
  reg [15:0] _T_157_0; 
  reg [31:0] _RAND_157;

  reg [15:0] _T_164_0; 
  reg [31:0] _RAND_164;
  reg [15:0] _T_165_0;
  reg [31:0] _RAND_165;
  reg [15:0] _T_166_0;
  reg [31:0] _RAND_166;
  reg [15:0] _T_167_0;
  reg [31:0] _RAND_167;

  reg [15:0] _T_174_0; 
  reg [31:0] _RAND_174;
  reg [15:0] _T_175_0;
  reg [31:0] _RAND_175;
  reg [15:0] _T_176_0;
  reg [31:0] _RAND_176;
  reg [15:0] _T_177_0;
  reg [31:0] _RAND_177;

  reg [15:0] _T_184_0; 
  reg [31:0] _RAND_184;
  reg [15:0] _T_185_0;
  reg [31:0] _RAND_185;
  reg [15:0] _T_186_0;
  reg [31:0] _RAND_186;
  reg [15:0] _T_187_0;
  reg [31:0] _RAND_187;
  

  reg  _T_236; 
  reg [31:0] _RAND_236;
  reg  _T_239; 
  reg [31:0] _RAND_238;
  reg  _T_242; 
  reg [31:0] _RAND_240;
  reg  _T_245; 
  reg [31:0] _RAND_242;
  

  reg  _T_262; 
  reg [31:0] _RAND_255;
  reg  _T_265; 
  reg [31:0] _RAND_257;
  reg  _T_268; 
  reg [31:0] _RAND_259;
  reg  _T_271; 
  reg [31:0] _RAND_261;

  reg  _T_288; 
  reg [31:0] _RAND_274;
  reg  _T_291; 
  reg [31:0] _RAND_276;
  reg  _T_294; 
  reg [31:0] _RAND_278;
  reg  _T_297; 
  reg [31:0] _RAND_280;
  

  reg  _T_314; 
  reg [31:0] _RAND_293;
  reg  _T_317; 
  reg [31:0] _RAND_295;
  reg  _T_320; 
  reg [31:0] _RAND_297;
  reg  _T_323; 
  reg [31:0] _RAND_299;
  
  
  
  
  
  //Tile/PE Instances
  Tile mesh_0_0 ( 
    .clock(mesh_0_0_clock),
    .io_in_a_0(mesh_0_0_io_in_a_0),
    .io_in_b_0(mesh_0_0_io_in_b_0),
    .io_in_d_0(mesh_0_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate),
    .io_out_a_0(mesh_0_0_io_out_a_0),
    .io_out_c_0(mesh_0_0_io_out_c_0),
    .io_out_b_0(mesh_0_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_0_io_out_control_0_propagate)
  );
  Tile mesh_0_1 ( 
    .clock(mesh_0_1_clock),
    .io_in_a_0(mesh_0_1_io_in_a_0),
    .io_in_b_0(mesh_0_1_io_in_b_0),
    .io_in_d_0(mesh_0_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate),
    .io_out_a_0(mesh_0_1_io_out_a_0),
    .io_out_c_0(mesh_0_1_io_out_c_0),
    .io_out_b_0(mesh_0_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_1_io_out_control_0_propagate)
  );
  Tile mesh_0_2 ( 
    .clock(mesh_0_2_clock),
    .io_in_a_0(mesh_0_2_io_in_a_0),
    .io_in_b_0(mesh_0_2_io_in_b_0),
    .io_in_d_0(mesh_0_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate),
    .io_out_a_0(mesh_0_2_io_out_a_0),
    .io_out_c_0(mesh_0_2_io_out_c_0),
    .io_out_b_0(mesh_0_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_2_io_out_control_0_propagate)
  );
  Tile mesh_0_3 (
    .clock(mesh_0_3_clock),
    .io_in_a_0(mesh_0_3_io_in_a_0),
    .io_in_b_0(mesh_0_3_io_in_b_0),
    .io_in_d_0(mesh_0_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate),
    .io_out_a_0(mesh_0_3_io_out_a_0),
    .io_out_c_0(mesh_0_3_io_out_c_0),
    .io_out_b_0(mesh_0_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_3_io_out_control_0_propagate)
  );
   Tile mesh_1_0 ( 
    .clock(mesh_1_0_clock),
    .io_in_a_0(mesh_1_0_io_in_a_0),
    .io_in_b_0(mesh_1_0_io_in_b_0),
    .io_in_d_0(mesh_1_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate),
    .io_out_a_0(mesh_1_0_io_out_a_0),
    .io_out_c_0(mesh_1_0_io_out_c_0),
    .io_out_b_0(mesh_1_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_0_io_out_control_0_propagate)
  );
  Tile mesh_1_1 ( 
    .clock(mesh_1_1_clock),
    .io_in_a_0(mesh_1_1_io_in_a_0),
    .io_in_b_0(mesh_1_1_io_in_b_0),
    .io_in_d_0(mesh_1_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate),
    .io_out_a_0(mesh_1_1_io_out_a_0),
    .io_out_c_0(mesh_1_1_io_out_c_0),
    .io_out_b_0(mesh_1_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_1_io_out_control_0_propagate)
     );
  Tile mesh_1_2 ( 
    .clock(mesh_1_2_clock),
    .io_in_a_0(mesh_1_2_io_in_a_0),
    .io_in_b_0(mesh_1_2_io_in_b_0),
    .io_in_d_0(mesh_1_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate),
    .io_out_a_0(mesh_1_2_io_out_a_0),
    .io_out_c_0(mesh_1_2_io_out_c_0),
    .io_out_b_0(mesh_1_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_2_io_out_control_0_propagate)
      );
  Tile mesh_1_3 ( 
    .clock(mesh_1_3_clock),
    .io_in_a_0(mesh_1_3_io_in_a_0),
    .io_in_b_0(mesh_1_3_io_in_b_0),
    .io_in_d_0(mesh_1_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate),
    .io_out_a_0(mesh_1_3_io_out_a_0),
    .io_out_c_0(mesh_1_3_io_out_c_0),
    .io_out_b_0(mesh_1_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_3_io_out_control_0_propagate)
      );
   Tile mesh_2_0 ( 
    .clock(mesh_2_0_clock),
    .io_in_a_0(mesh_2_0_io_in_a_0),
    .io_in_b_0(mesh_2_0_io_in_b_0),
    .io_in_d_0(mesh_2_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate),
    .io_out_a_0(mesh_2_0_io_out_a_0),
    .io_out_c_0(mesh_2_0_io_out_c_0),
    .io_out_b_0(mesh_2_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_0_io_out_control_0_propagate)
     );
  Tile mesh_2_1 ( 
    .clock(mesh_2_1_clock),
    .io_in_a_0(mesh_2_1_io_in_a_0),
    .io_in_b_0(mesh_2_1_io_in_b_0),
    .io_in_d_0(mesh_2_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate),
    .io_out_a_0(mesh_2_1_io_out_a_0),
    .io_out_c_0(mesh_2_1_io_out_c_0),
    .io_out_b_0(mesh_2_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_1_io_out_control_0_propagate)
     );
  Tile mesh_2_2 (
    .clock(mesh_2_2_clock),
    .io_in_a_0(mesh_2_2_io_in_a_0),
    .io_in_b_0(mesh_2_2_io_in_b_0),
    .io_in_d_0(mesh_2_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate),
    .io_out_a_0(mesh_2_2_io_out_a_0),
    .io_out_c_0(mesh_2_2_io_out_c_0),
    .io_out_b_0(mesh_2_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_2_io_out_control_0_propagate)
     );
  Tile mesh_2_3 ( 
    .clock(mesh_2_3_clock),
    .io_in_a_0(mesh_2_3_io_in_a_0),
    .io_in_b_0(mesh_2_3_io_in_b_0),
    .io_in_d_0(mesh_2_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate),
    .io_out_a_0(mesh_2_3_io_out_a_0),
    .io_out_c_0(mesh_2_3_io_out_c_0),
    .io_out_b_0(mesh_2_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_3_io_out_control_0_propagate)
     );
    Tile mesh_3_0 ( 
    .clock(mesh_3_0_clock),
    .io_in_a_0(mesh_3_0_io_in_a_0),
    .io_in_b_0(mesh_3_0_io_in_b_0),
    .io_in_d_0(mesh_3_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate),
    .io_out_a_0(mesh_3_0_io_out_a_0),
    .io_out_c_0(mesh_3_0_io_out_c_0),
    .io_out_b_0(mesh_3_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_0_io_out_control_0_propagate)
  );
  Tile mesh_3_1 ( 
    .clock(mesh_3_1_clock),
    .io_in_a_0(mesh_3_1_io_in_a_0),
    .io_in_b_0(mesh_3_1_io_in_b_0),
    .io_in_d_0(mesh_3_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate),
    .io_out_a_0(mesh_3_1_io_out_a_0),
    .io_out_c_0(mesh_3_1_io_out_c_0),
    .io_out_b_0(mesh_3_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_1_io_out_control_0_propagate)
  );
  Tile mesh_3_2 ( 
    .clock(mesh_3_2_clock),
    .io_in_a_0(mesh_3_2_io_in_a_0),
    .io_in_b_0(mesh_3_2_io_in_b_0),
    .io_in_d_0(mesh_3_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate),
    .io_out_a_0(mesh_3_2_io_out_a_0),
    .io_out_c_0(mesh_3_2_io_out_c_0),
    .io_out_b_0(mesh_3_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_2_io_out_control_0_propagate)
  );
  Tile mesh_3_3 ( 
    .clock(mesh_3_3_clock),
    .io_in_a_0(mesh_3_3_io_in_a_0),
    .io_in_b_0(mesh_3_3_io_in_b_0),
    .io_in_d_0(mesh_3_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate),
    .io_out_a_0(mesh_3_3_io_out_a_0),
    .io_out_c_0(mesh_3_3_io_out_c_0),
    .io_out_b_0(mesh_3_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_3_io_out_control_0_propagate)
   );
   
//Final Ouput Register at Bottom  
always @(posedge clock) begin
  io_out_c_0_0 <= mesh_3_0_io_out_c_0; 
  io_out_c_1_0 <= mesh_3_1_io_out_c_0; 
  io_out_c_2_0 <= mesh_3_2_io_out_c_0; 
  io_out_c_3_0 <= mesh_3_3_io_out_c_0; 
end

 //Mesh Internal input/ouput wires Connections
  assign mesh_0_0_clock = clock; 	  
  assign mesh_0_0_io_in_a_0 = _T_1_0; 
  assign mesh_0_0_io_in_b_0 = _T_74_0;
  assign mesh_0_0_io_in_d_0 = _T_154_0; 
  assign mesh_0_0_io_in_control_0_propagate = _T_236; 
  
  assign mesh_0_1_clock = clock; 		
  assign mesh_0_1_io_in_a_0 = _T_2_0; 	
  assign mesh_0_1_io_in_b_0 = _T_84_0; 
  assign mesh_0_1_io_in_d_0 = _T_164_0;
  assign mesh_0_1_io_in_control_0_propagate = _T_262; 
  
  assign mesh_0_2_clock = clock; 		
  assign mesh_0_2_io_in_a_0 = _T_3_0; 	
  assign mesh_0_2_io_in_b_0 = _T_94_0; 
  assign mesh_0_2_io_in_d_0 = _T_174_0;
  assign mesh_0_2_io_in_control_0_propagate = _T_288; 
  
  assign mesh_0_3_clock = clock; 		
  assign mesh_0_3_io_in_a_0 = _T_4_0; 	
  assign mesh_0_3_io_in_b_0 = _T_104_0;
  assign mesh_0_3_io_in_d_0 = _T_184_0;
  assign mesh_0_3_io_in_control_0_propagate = _T_314; 
  
  assign mesh_1_0_clock = clock; 		
  assign mesh_1_0_io_in_a_0 = _T_10_0; 	
  assign mesh_1_0_io_in_b_0 = _T_75_0; 	
  assign mesh_1_0_io_in_d_0 = _T_155_0; 
  assign mesh_1_0_io_in_control_0_propagate = _T_239; 
  assign mesh_1_1_clock = clock; 		
  assign mesh_1_1_io_in_a_0 = _T_11_0; 
  assign mesh_1_1_io_in_b_0 = _T_85_0; 
  assign mesh_1_1_io_in_d_0 = _T_165_0;
  assign mesh_1_1_io_in_control_0_propagate = _T_265; 
  assign mesh_1_2_clock = clock; 		
  assign mesh_1_2_io_in_a_0 = _T_12_0; 
  assign mesh_1_2_io_in_b_0 = _T_95_0; 
  assign mesh_1_2_io_in_d_0 = _T_175_0;
  assign mesh_1_2_io_in_control_0_propagate = _T_291; 
  assign mesh_1_3_clock = clock; 		
  assign mesh_1_3_io_in_a_0 = _T_13_0; 
  assign mesh_1_3_io_in_b_0 = _T_105_0;
  assign mesh_1_3_io_in_d_0 = _T_185_0;
  assign mesh_1_3_io_in_control_0_propagate = _T_317; 
  
  assign mesh_2_0_clock = clock; 		
  assign mesh_2_0_io_in_a_0 = _T_19_0; 
  assign mesh_2_0_io_in_b_0 = _T_76_0; 
  assign mesh_2_0_io_in_d_0 = _T_156_0;
  assign mesh_2_0_io_in_control_0_propagate = _T_242; 
  assign mesh_2_1_clock = clock; 		
  assign mesh_2_1_io_in_a_0 = _T_20_0; 
  assign mesh_2_1_io_in_b_0 = _T_86_0; 
  assign mesh_2_1_io_in_d_0 = _T_166_0;
  assign mesh_2_1_io_in_control_0_propagate = _T_268; 
  assign mesh_2_2_clock = clock; 		
  assign mesh_2_2_io_in_a_0 = _T_21_0; 
  assign mesh_2_2_io_in_b_0 = _T_96_0; 
  assign mesh_2_2_io_in_d_0 = _T_176_0;
  assign mesh_2_2_io_in_control_0_propagate = _T_294; 
  assign mesh_2_3_clock = clock; 		
  assign mesh_2_3_io_in_a_0 = _T_22_0; 
  assign mesh_2_3_io_in_b_0 = _T_106_0;
  assign mesh_2_3_io_in_d_0 = _T_186_0;
  assign mesh_2_3_io_in_control_0_propagate = _T_320; 
  
  assign mesh_3_0_clock = clock; 		
  assign mesh_3_0_io_in_a_0 = _T_28_0; 
  assign mesh_3_0_io_in_b_0 = _T_77_0; 
  assign mesh_3_0_io_in_d_0 = _T_157_0;
  assign mesh_3_0_io_in_control_0_propagate = _T_245; 
  assign mesh_3_1_clock = clock; 		
  assign mesh_3_1_io_in_a_0 = _T_29_0; 
  assign mesh_3_1_io_in_b_0 = _T_87_0; 
  assign mesh_3_1_io_in_d_0 = _T_167_0;
  assign mesh_3_1_io_in_control_0_propagate = _T_271; 
  assign mesh_3_2_clock = clock; 		
  assign mesh_3_2_io_in_a_0 = _T_30_0; 
  assign mesh_3_2_io_in_b_0 = _T_97_0; 
  assign mesh_3_2_io_in_d_0 = _T_177_0;
  assign mesh_3_2_io_in_control_0_propagate = _T_297; 
  assign mesh_3_3_clock = clock; 		
  assign mesh_3_3_io_in_a_0 = _T_31_0; 
  assign mesh_3_3_io_in_b_0 = _T_107_0;
  assign mesh_3_3_io_in_d_0 = _T_187_0;
  assign mesh_3_3_io_in_control_0_propagate = _T_323; 
  
//Random values to assign registers  
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4_0 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
 
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10_0 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11_0 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12_0 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13_0 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19_0 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20_0 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21_0 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22_0 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
 
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_28_0 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29_0 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30_0 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_31_0 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  

  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_74_0 = _RAND_74[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_75_0 = _RAND_75[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_76_0 = _RAND_76[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77_0 = _RAND_77[7:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_84_0 = _RAND_84[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_85_0 = _RAND_85[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_86_0 = _RAND_86[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_87_0 = _RAND_87[7:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_94_0 = _RAND_94[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_95_0 = _RAND_95[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_96_0 = _RAND_96[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_97_0 = _RAND_97[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_98_0 = _RAND_98[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_99_0 = _RAND_99[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_100_0 = _RAND_100[7:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_101_0 = _RAND_101[7:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_104_0 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_105_0 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_106_0 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_107_0 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_154_0 = _RAND_154[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_155_0 = _RAND_155[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_156_0 = _RAND_156[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_157_0 = _RAND_157[15:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_164_0 = _RAND_164[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_165_0 = _RAND_165[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_166_0 = _RAND_166[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_167_0 = _RAND_167[15:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_174_0 = _RAND_174[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_175_0 = _RAND_175[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_176_0 = _RAND_176[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_177_0 = _RAND_177[15:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_184_0 = _RAND_184[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_185_0 = _RAND_185[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_186_0 = _RAND_186[15:0] ;
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_187_0 = _RAND_187[15:0] ;
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_236 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_239 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_242 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_245 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_262 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_265 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_268 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_271 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT

  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_288 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_291 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_294 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_297 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_314 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_317 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_320 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_323 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
  //A input Registers conenction for column 0
    _T_1_0 <= io_in_a_0_0;
    _T_2_0 <= mesh_0_0_io_out_a_0;
    _T_3_0 <= mesh_0_1_io_out_a_0;
    _T_4_0 <= mesh_0_2_io_out_a_0;
	
  //A input Registers conenction for column 1
    _T_10_0 <= io_in_a_1_0;
    _T_11_0 <= mesh_1_0_io_out_a_0;
    _T_12_0 <= mesh_1_1_io_out_a_0;
    _T_13_0 <= mesh_1_2_io_out_a_0;

//A input Registers conenction for column 2
    _T_19_0 <= io_in_a_2_0;
    _T_20_0 <= mesh_2_0_io_out_a_0;
    _T_21_0 <= mesh_2_1_io_out_a_0;
    _T_22_0 <= mesh_2_2_io_out_a_0;

//A input Registers conenction for column 3
    _T_28_0 <= io_in_a_3_0;;
    _T_29_0 <= mesh_3_0_io_out_a_0;
    _T_30_0 <= mesh_3_1_io_out_a_0;
    _T_31_0 <= mesh_3_2_io_out_a_0;


    _T_74_0 <= io_in_d_0_0;
    _T_75_0 <= mesh_0_0_io_out_b_0;
    _T_76_0 <= mesh_1_0_io_out_b_0;
    _T_77_0 <= mesh_2_0_io_out_b_0;
 
    _T_84_0 <= io_in_d_1_0;
    _T_85_0 <= mesh_0_1_io_out_b_0;
    _T_86_0 <= mesh_1_1_io_out_b_0;
    _T_87_0 <= mesh_2_1_io_out_b_0;
    

    _T_94_0 <=  io_in_d_2_0;
    _T_95_0 <= mesh_0_2_io_out_b_0;
    _T_96_0 <= mesh_1_2_io_out_b_0;
    _T_97_0 <= mesh_2_2_io_out_b_0;
    

    _T_104_0 <= io_in_d_3_0;
    _T_105_0 <= mesh_0_3_io_out_b_0;
    _T_106_0 <= mesh_1_3_io_out_b_0;
    _T_107_0 <= mesh_2_3_io_out_b_0;
 
    _T_154_0 <= io_in_b_0_0;
    _T_155_0 <= mesh_0_0_io_out_c_0;
    _T_156_0 <= mesh_1_0_io_out_c_0;
    _T_157_0 <= mesh_2_0_io_out_c_0;
    

    _T_164_0 <= io_in_b_1_0;
    _T_165_0 <= mesh_0_1_io_out_c_0;
    _T_166_0 <= mesh_1_1_io_out_c_0;
    _T_167_0 <= mesh_2_1_io_out_c_0;
    

    _T_174_0 <= io_in_b_2_0;
    _T_175_0 <= mesh_0_2_io_out_c_0;
    _T_176_0 <= mesh_1_2_io_out_c_0;
    _T_177_0 <= mesh_2_2_io_out_c_0;
    
	
    _T_184_0 <= io_in_b_3_0;
    _T_185_0 <= mesh_0_3_io_out_c_0;
    _T_186_0 <= mesh_1_3_io_out_c_0;
    _T_187_0 <= mesh_2_3_io_out_c_0;
    
//CTL_PROP input Registers conenction for column 0	
    _T_236 <= io_in_control_0_0_propagate;
    _T_239 <= mesh_0_0_io_out_control_0_propagate;
    _T_242 <= mesh_1_0_io_out_control_0_propagate;
    _T_245 <= mesh_2_0_io_out_control_0_propagate;
    
//CTL_PROP input Registers conenction for column 1
	_T_262 <=io_in_control_1_0_propagate;
    _T_265 <= mesh_0_1_io_out_control_0_propagate;
    _T_268 <= mesh_1_1_io_out_control_0_propagate;
    _T_271 <= mesh_2_1_io_out_control_0_propagate;
    
//CTL_PROP input Registers conenction for column 2
    _T_288 <=  io_in_control_2_0_propagate;
    _T_291 <= mesh_0_2_io_out_control_0_propagate;
    _T_294 <= mesh_1_2_io_out_control_0_propagate;
    _T_297 <= mesh_2_2_io_out_control_0_propagate;
    
//CTL_PROP input Registers conenction for column 3	
    _T_314 <= io_in_control_3_0_propagate;
    _T_317 <= mesh_0_3_io_out_control_0_propagate;
    _T_320 <= mesh_1_3_io_out_control_0_propagate;
    _T_323 <= mesh_2_3_io_out_control_0_propagate;
    
	
  end
endmodule
